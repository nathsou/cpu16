module ROM (
    input logic [15:0] addr,
    output logic [15:0] data
);
    always_comb begin
        case (addr)
            16'h0000: data = 16'h71FF;
            16'h0001: data = 16'h48BA;
            16'h0002: data = 16'h6808;
            16'h0003: data = 16'hC9BA;
            16'h0004: data = 16'h68BA;
            16'h0005: data = 16'hC9B8;
            16'h0006: data = 16'h5020;
            16'h0007: data = 16'h6805;
            16'h0008: data = 16'hEDE0;
            16'h0009: data = 16'hAE00;
            16'h000A: data = 16'hF614;
            16'h000B: data = 16'h680A;
            16'h000C: data = 16'hFFA0;
            16'h000D: data = 16'h4820;
            16'h000E: data = 16'h5000;
            16'h000F: data = 16'h6805;
            16'h0010: data = 16'hEDE0;
            16'h0011: data = 16'hAE00;
            16'h0012: data = 16'hF614;
            16'h0013: data = 16'h6846;
            16'h0014: data = 16'hFFA0;
            16'h0015: data = 16'h0000;
            16'h0016: data = 16'h8800;
            16'h0017: data = 16'h9001;
            16'h0018: data = 16'h4802;
            16'h0019: data = 16'h5027;
            16'h001A: data = 16'h6808;
            16'h001B: data = 16'hD2BA;
            16'h001C: data = 16'h6810;
            16'h001D: data = 16'hD2B8;
            16'h001E: data = 16'h9100;
            16'h001F: data = 16'h53E8;
            16'h0020: data = 16'h9101;
            16'h0021: data = 16'h5064;
            16'h0022: data = 16'h9102;
            16'h0023: data = 16'h500A;
            16'h0024: data = 16'h9103;
            16'h0025: data = 16'h5001;
            16'h0026: data = 16'h9104;
            16'h0027: data = 16'h8882;
            16'h0028: data = 16'h8880;
            16'h0029: data = 16'hC101;
            16'h002A: data = 16'h6807;
            16'h002B: data = 16'hFFA8;
            16'h002C: data = 16'h9081;
            16'h002D: data = 16'h6830;
            16'h002E: data = 16'hAA00;
            16'h002F: data = 16'h8201;
            16'h0030: data = 16'hF615;
            16'h0031: data = 16'hBE80;
            16'h0032: data = 16'h4800;
            16'h0033: data = 16'h5000;
            16'h0034: data = 16'h6805;
            16'h0035: data = 16'hC1A1;
            16'h0036: data = 16'h681E;
            16'h0037: data = 16'hFFA4;
            16'h0038: data = 16'h6000;
            16'h0039: data = 16'h9982;
            16'h003A: data = 16'hA880;
            16'h003B: data = 16'hC561;
            16'h003C: data = 16'h6807;
            16'h003D: data = 16'hFFB0;
            16'h003E: data = 16'hA880;
            16'h003F: data = 16'hED61;
            16'h0040: data = 16'hA800;
            16'h0041: data = 16'hE414;
            16'h0042: data = 16'h680A;
            16'h0043: data = 16'hFFA1;
            16'h0044: data = 16'hC914;
            16'h0045: data = 16'hC040;
            16'h0046: data = 16'h6806;
            16'h0047: data = 16'hFFA8;
            16'h0048: data = 16'hC080;
            16'h0049: data = 16'h6803;
            16'h004A: data = 16'hFFA8;
            16'h004B: data = 16'h6818;
            16'h004C: data = 16'hFFA1;
            16'h004D: data = 16'h9881;
            16'h004E: data = 16'hDB40;
            16'h004F: data = 16'h6830;
            16'h0050: data = 16'hED80;
            16'h0051: data = 16'hAB00;
            16'h0052: data = 16'hD214;
            16'h0053: data = 16'h6820;
            16'h0054: data = 16'hFFA1;
            16'h0055: data = 16'h8881;
            16'h0056: data = 16'hC940;
            16'h0057: data = 16'h8100;
            16'h0058: data = 16'hF615;
            16'h0059: data = 16'hBE80;
            16'h005A: data = 16'h6000;
            16'h005B: data = 16'hE415;
            16'h005C: data = 16'h9980;
            16'h005D: data = 16'h9864;
            16'h005E: data = 16'hC301;
            16'h005F: data = 16'h680D;
            16'h0060: data = 16'hFFA4;
            16'h0061: data = 16'h5880;
            16'h0062: data = 16'h6808;
            16'h0063: data = 16'hDBBA;
            16'h0064: data = 16'hDB18;
            16'h0065: data = 16'hDB40;
            16'h0066: data = 16'h9C00;
            16'h0067: data = 16'hD214;
            16'h0068: data = 16'h98E4;
            16'h0069: data = 16'h9C00;
            16'h006A: data = 16'hC914;
            16'h006B: data = 16'h6810;
            16'h006C: data = 16'hFFA1;
            16'h006D: data = 16'hF615;
            16'h006E: data = 16'hBE80;
            default: data = 16'h0000;
        endcase
    end
endmodule
