module veryl_Top;
    initial begin
        $display("Hello, world!");
    end
endmodule
//# sourceMappingURL=Top.sv.map
